C00|Lip_Proper
C01|Root_Of_Tongue
C02|Root_Of_Tongue
C03|Sublingual_Region
C07|Salivary_Gland
C09|Pharynx
C11|Posterior_Wall_Of_The_Nasopharynx
C12|Hypopharynx
C14|Pharynx
C15|Esophagus
C16|Stomach
C17|Small_Intestine
C18|Appendix
C20|Rectal
C21|Anal_Canal
C22|Intrahepatic_Bile_Duct
C23|Extrahepatic_Bile_Duct
C25|Pancreas
C26|Entire_Digestive_Organ
C30|Middle_Ear
C31|Nasal_Sinus
C32|Larynx
C33|Trachea
C34|Bronchus
C37|Thymus_Gland
C38|Pleura
C39|Respiratory_System
C40|Mandible
C41|Mandible
C42|Reticuloendothelial_System
C44|Skin
C47|Peripheral_Nerve
C48|Retroperitoneal_Space
C50|Breast
C51|Vulva
C53|Cervix_Uteri
C54|Corpus_Uteri
C55|Uterus
C56|Ovary
C57|Fallopian_Tube
C58|Placenta_Part
C60|Penis
C61|Prostate
C62|Testis
C63|Scrotum
C64|Kidney
C65|Renal_Pelvis
C67|Urinary_Bladder
C68|Genitourinary_System
C69|Eye
C70|Meninges
C71|Cerebellum
C72|Central_Nervous_System
C73|Thyroid_Gland
C74|Adrenal_Gland
C75|Endocrine_Gland
C77|Lymph_Node
C80|Undetermined
